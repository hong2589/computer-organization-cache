`include "opcodes.v"
`define WORD_SIZE 16    // data and address word size
module cache(

);
endmodule